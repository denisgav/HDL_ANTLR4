﻿entity some_test_bench is
end some_test_bench;

architecture some_test_bench of some_test_bench is
	subtype  my_real is real range 0.0 to 1024.0; 
	subtype natural is integer range 0 to integer'high; 
	subtype positive is integer range 1 to integer'high; 
begin
end architecture some_test_bench;