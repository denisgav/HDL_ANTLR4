entity some_test_bench is
end entity;

architecture some_test_bench of some_test_bench is
	signal x1, x2, x3, x4 : bit;
	signal y1, y2, y3, y4 : bit;
begin


end architecture some_test_bench;